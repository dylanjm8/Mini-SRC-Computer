// DIV datapath_tb.v file: <This is the filename>
`timescale 1ns/10ps
module div_tb();
	reg PCout,Zlowout, Zhighout, MDRout, R2out, R3out; // add any other signals to see in your simulation
	reg MARin, Zin, PCin, MDRin, IRin, Yin, LOin, HIin;
	reg IncPC, Read, DIV, R1in, R2in, R3in;
	reg Clock;
	reg [31:0] Mdatain;
	reg clear;
	
	
Datapath DUT(PCout, Zlowout, Zhighout, MDRout, R2out, R3out, MARin, Zin, PCin, MDRin, IRin, Yin, LOin, HIin, IncPC, Read, DIV, R1in,
R2in, R3in, Clock, Mdatain, clear);

	 parameter Default = 4'b0000, Reg_load1= 4'b0001, Reg_load1b= 4'b0010,
					Reg_load2= 4'b0011, Reg_load2b = 4'b0100, Reg_load3 = 4'b0101,
					Reg_load3b = 4'b0110, T0= 4'b0111, T1= 4'b1000,T2= 4'b1001, T3= 4'b1010, T4= 4'b1011, T5= 4'b1100, T6= 4'b1101;
	reg [3:0] Present_state = Default;
// add test logic here
initial
	begin
	Clock = 0;
	forever #10 Clock = ~ Clock;
end

always @(posedge Clock) // finite state machine; if clock rising-edge
	begin
		case (Present_state)
			Default : Present_state = Reg_load1;
			Reg_load1 : Present_state = Reg_load1b;
			Reg_load1b : Present_state = Reg_load2;
			Reg_load2 : Present_state = Reg_load2b;
			Reg_load2b : Present_state = Reg_load3;
			Reg_load3 : Present_state = Reg_load3b;
			Reg_load3b : Present_state = T0;
			T0 : Present_state = T1;
			T1 : Present_state = T2;
			T2 : Present_state = T3;
			T3 : Present_state = T4;
			T4 : Present_state = T5;
			T5 : Present_state = T6;


		endcase
	end

always @(Present_state) // do the required job in each state
	begin
		case (Present_state) // assert the required signals in each clock cycle
			Default: begin
					clear <= 0; PCout <= 0; Zlowout <= 0; Zhighout <= 0; MDRout <= 0; // initialize the signals
					R2out <= 0; R3out <= 0; MARin <= 0; Zin <= 0;
					PCin <=0; MDRin <= 0; IRin <= 0; Yin <= 0; LOin <= 0; HIin <= 0;
					IncPC <= 0; Read <= 0; DIV <= 0;
					R1in <= 0; R2in <= 0; R3in <= 0; Mdatain <= 32'h00000000;
			end
			Reg_load1: begin
					Mdatain <= 32'h00000007;
					Read = 0; MDRin = 0; // the first zero is there for completeness
					MDRin <= 1; Read <= 1;
					#15 MDRin <= 0; Read <= 0;// implementation; same goes for the other states
			end
			Reg_load1b: begin
				 MDRout <= 1; R2in <= 1;
				#15 MDRout <= 0; R2in <= 0; // initialize R2 with the value $22
			end
			Reg_load2: begin
				Mdatain <= 32'h00000003;
				 Read <= 1; MDRin <= 1;
				#15 Read <= 0; MDRin <= 0;
			end
			Reg_load2b: begin
				 MDRout <= 1; R3in <= 1;
				#15 MDRout <= 0; R3in <= 0; // initialize R3 with the value $24
			end
			Reg_load3: begin
				Mdatain <= 32'h00000027;
				Read <= 1; MDRin <= 1;
				#15 Read <= 0; MDRin <= 0;
			end
			Reg_load3b: begin
				MDRout <= 1; R1in <= 1;
				#15 MDRout <= 0; R1in <= 0; // initialize R1 with the value $26
			end
		T0: begin // see if you need to de-assert these signals
			PCout <= 1; MARin <= 1; Zin <= 1;
		end
		T1: begin
			PCout <= 0; MARin <= 0; Zin <= 0;
			Zlowout <= 1; PCin <= 1; Read <= 1; MDRin <= 1; IncPC <= 1;
			Mdatain <= 32'h19180000; // opcode for “DIV R2, R3”

		end
		T2: begin
			Zlowout <= 0; PCin <= 0; Read <= 0; MDRin <= 0; IncPC <= 0;
			MDRout <= 1; IRin <= 1;
		end
		T3: begin
			MDRout <= 0; IRin <= 0;		
			R2out <= 1; Yin <= 1;
		end
		T4: begin
			R2out <= 0; Yin <= 0;
			R3out <= 1; DIV <= 1; Zin <= 1;
		end
		T5: begin
			R3out <= 0; DIV <= 0; Zin <= 0;
			Zlowout <= 1; LOin <= 1;
		end
		T6: begin
			Zlowout <= 0; LOin <= 0;
			Zhighout <= 1; HIin <= 1;
			#20 Zhighout <= 0; HIin <= 0; 
		end
	  endcase
	end
endmodule